//Testbench: ISSUE_QUEUE_MULT

`timescale 1ns / 100ps

module testbench;


endmodule
