//-----------------------------------------------------
// Design Name 	: RST
// File Name   	: rst.v
// Function    	: 
// Coder  	: 
// Other	:
//-----------------------------------------------------

module rst (
  	input        	clock,
  	input        	reset,

  	input  	[ 4:0] 	Rsaddr_rst,
  	output 	[ 4:0] 	Rstag_rst,
  	output       	Rsvalid_rst,

  	input  	[ 4:0] 	Rtaddr_rst,
  	output 	[ 4:0] 	Rttag_rst,
  	output       	Rtvalid_rst,
  
  	input  	[ 4:0] 	RB_tag_rst,
	input        	RB_valid_rst,

 	input  	[ 4:0] 	Wdata_rst,
  	input  	[ 4:0] 	Waddr_rst,
	input 	[31:0] 	Wen0_rst,
	input 		Wen_rst,
	output reg [31:0] 	Wen1_rst 
	);

reg 	[ 5:0] 	RST_reg 	[31:0];

wire 	[ 5:0]	CDB_Token;
reg 	[31:0]	Comparator;

integer i;
integer j;
integer k;
integer l;

always@(posedge clock or posedge reset) begin
	if(reset) begin
		for (i=0; i < 32; i=i+1 ) begin
      			RST_reg [i] <= 6'b0_00000; //se ponen todos los registros como no validos.
			Wen1_rst[i] <= 0;
		end
    	end else begin   
      		if(Wen_rst) begin
        		RST_reg [Waddr_rst] <= {1'b1, Wdata_rst};
      		end 
     /*  falta borrar los tags */
		if(|Wen0_rst) begin
			for (l=0; l < 32; l=l+1 ) begin
				if (Wen0_rst[l]) begin
        				RST_reg [l] <= {1'b0, 5'b0};
				end	
			end
		end 
    	end
end

always @* begin
	for (j=0; j< 32;j=j+1) begin
	 	Comparator [j] = (RST_reg[j] ~^ CDB_Token);
	end
end 

always @* begin
	for (k=0; k< 32;k=k+1) begin
	 	Wen1_rst [k] = Comparator[k] & (~Wen0_rst[k]);
	end
end 

assign CDB_Token = {RB_valid_rst,RB_tag_rst};

// Read Rs and Rt
assign Rstag_rst 	= RST_reg[Rsaddr_rst][4:0];
assign Rttag_rst 	= RST_reg[Rtaddr_rst][4:0];
assign Rsvalid_rst 	= RST_reg[Rsaddr_rst][  5];
assign Rtvalid_rst 	= RST_reg[Rtaddr_rst][  5];

endmodule
