//Testbench: ROB

`timescale 1ns / 100ps

module testbench;


endmodule
