//Testbench: Order_Queue_Mem

`timescale 1ns / 100ps

module testbench;


endmodule
