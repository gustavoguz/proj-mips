//Testbench: FULL_ADDER

`timescale 1ns / 100ps

module testbench;


endmodule
