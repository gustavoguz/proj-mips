
module tb_BackEnd();
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  
  


endmodule
