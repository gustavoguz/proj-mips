//Testbench: Coder32_5

`timescale 1ns / 100ps

module testbench;


endmodule
