//Testbench: RTS

`timescale 1ns / 100ps

module testbench;


endmodule
