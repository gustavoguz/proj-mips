//Testbench: ISSUE_QUEUE_INT

`timescale 1ns / 100ps

module testbench;


endmodule
