//Testbench: XOR

`timescale 1ns / 100ps

module testbench;


endmodule
