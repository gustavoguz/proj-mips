//Testbench: ADDRESS_LOGIC

`timescale 1ns / 100ps

module testbench;


endmodule
