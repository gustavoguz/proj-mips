//Testbench: FULL_ADDER_32

`timescale 1ns / 100ps

module testbench;


endmodule
