//Testbench: ISSUE_UNIT

`timescale 1ns / 100ps

module testbench;


endmodule
