//Testbench: RAM

`timescale 1ns / 100ps

module testbench;


endmodule
