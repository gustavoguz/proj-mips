//Testbench: ISSUE_QUEUE_LS

`timescale 1ns / 100ps

module testbench;


endmodule
